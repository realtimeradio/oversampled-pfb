`timescale 1ns / 1ps
`default_nettype none

module symbolicpe (
  input wire logic clk,
  input string din,
  input string coeff,
  input string sin,
  output string sout
);

endmodule
